
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07/26/2025 02:05:08 PM
// Design Name: 
// Module Name: fifo2axis
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module fifo2axis #(
    parameter DATA_WIDTH = 32,
    parameter THRESHOLD = 4,
    parameter DEPTH = 10
)(
    input  wire        clk,
    input  wire        rst,

    // FIFO interface
    input  wire [31:0] fifo_data,
    input  wire        data_ready,

    // AXI Stream master
    output reg [31:0]  s_axis_tdata,
    output reg         s_axis_tvalid,
    input  wire        s_axis_tready,
    output wire        start_hls,
    input wire         s_axis_tlast
);

    // States
    localparam IDLE       = 3'd0,
               READ_FIFO  = 3'd1,
               WAIT_START = 3'd2,
               SEND       = 3'd3,
               DONE       = 3'd4;

    reg [2:0] state, next_state;

    // Internal buffer
    reg [31:0] buffer [0:3];
    reg [1:0]  buffer_index;
    reg [1:0]  send_index;
    reg start_hls_module;
    
    // When RESET signal is 0 and module starts, also start the HLS module
    assign start_hls = ~rst; 

    // FSM Sequential
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            state <= IDLE;
            buffer_index <= 2'd0;
            send_index <= 2'd0;
            s_axis_tvalid <= 0;
            s_axis_tdata  <= 32'd0;
            
        end else begin
            state = next_state;
            
            case (state)
                IDLE: begin
                    if (data_ready) begin
                        next_state <= READ_FIFO;
                    end else begin
                    	next_state <= IDLE;
                        buffer_index <= 0;
                    end
                end
               
                READ_FIFO: begin
                    buffer[buffer_index] <= fifo_data;
                    
                    if (buffer_index == 2'd3) begin
                        next_state <= WAIT_START;
                    end else begin
                        buffer_index <= buffer_index + 1;
                        next_state <= READ_FIFO;
                    end
                end

                WAIT_START: begin
                    if (s_axis_tready) begin
                        send_index <= 0;
                        next_state <= SEND;
                    end else begin
                        next_state <= WAIT_START;
                    end
                end
                
                SEND: begin
                    
                    #5; //wait a bit for AXISTREAM MODULE
                    
                    if (s_axis_tready) begin
                        s_axis_tdata  <= buffer[send_index];
                        s_axis_tvalid <= 1;
                        #10
                        s_axis_tvalid <= 0;
                        
                        if (send_index == 2'd3) begin
                            next_state = DONE;
                        end else begin
                            send_index <= send_index + 1;
                            next_state <= SEND;
                        end

                    end else begin
                        next_state <= SEND;
                    end

                end
                
                
                DONE: begin
                    if (s_axis_tlast) begin
                        s_axis_tdata = {32{1'bx}};
                        next_state <= IDLE;
                    end else begin
                        next_state <= DONE;
                    end
                end
                
                default: begin
                    next_state <= IDLE;
                end
            endcase
        end
    end

endmodule
